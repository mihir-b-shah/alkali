module ep2top#()
(
	 input  wire clk, 
	 input  wire rst,
	//input ports BUF
	input wire [512-1:0] NET_RECV_0_tdata ,
	input wire [64-1:0] NET_RECV_0_tkeep ,
	input wire  NET_RECV_0_tlast ,
	input wire  NET_RECV_0_tvalid ,
	output wire  NET_RECV_0_tready,
	//output ports BUF
	output wire [512-1:0] NET_SEND_0_tdata ,
	output wire [64-1:0] NET_SEND_0_tkeep ,
	output wire  NET_SEND_0_tlast ,
	output wire  NET_SEND_0_tvalid ,
	input wire  NET_SEND_0_tready
);
atom_CAM#(
)err_tracker_table_3(
	 .clk(clk), 
	 .rst(rst) ,
	//lookup port 
	.s_lookup_req_index({err_tracker_table_3lookup_p_0_req_index}),
	.s_lookup_req_valid({err_tracker_table_3lookup_p_0_req_valid}),
	.s_lookup_req_ready({err_tracker_table_3lookup_p_0_req_ready}),
	.s_lookup_value_valid({err_tracker_table_3lookup_p_0_value_valid}),
	.s_lookup_value_data({err_tracker_table_3lookup_p_0_value_data}),
	.s_lookup_value_ready({err_tracker_table_3lookup_p_0_value_ready}),
	//update port 
	.s_update_req_index({err_tracker_table_3update_p_0_req_index}),
	.s_update_req_index_valid({err_tracker_table_3update_p_0_req_index_valid}),
	.s_update_req_index_ready({err_tracker_table_3update_p_0_req_index_ready}),
	.s_update_req_data({err_tracker_table_3update_p_0_req_data}),
	.s_update_req_data_valid({err_tracker_table_3update_p_0_req_data_valid}),
	.s_update_req_data_ready({err_tracker_table_3update_p_0_req_data_ready})
);

//Table lookup port wire def 
 wire [32-1:0] err_tracker_table_3lookup_p_0_req_index;
 wire  err_tracker_table_3lookup_p_0_req_valid;
 wire  err_tracker_table_3lookup_p_0_req_ready;
 wire  err_tracker_table_3lookup_p_0_value_valid;
 wire  err_tracker_table_3lookup_p_0_value_ready;
 wire [96-1:0] err_tracker_table_3lookup_p_0_value_data;

//Table update port wire def 
 wire [32-1:0] err_tracker_table_3update_p_0_req_index;
 wire  err_tracker_table_3update_p_0_req_index_valid;
 wire  err_tracker_table_3update_p_0_req_index_ready;
 wire [96-1:0] err_tracker_table_3update_p_0_req_data;
 wire  err_tracker_table_3update_p_0_req_data_valid;
 wire  err_tracker_table_3update_p_0_req_data_ready;

atom_CAM#(
)firewall_tcpport_table_0(
	 .clk(clk), 
	 .rst(rst) ,
	//lookup port 
	.s_lookup_req_index({firewall_tcpport_table_0lookup_p_0_req_index}),
	.s_lookup_req_valid({firewall_tcpport_table_0lookup_p_0_req_valid}),
	.s_lookup_req_ready({firewall_tcpport_table_0lookup_p_0_req_ready}),
	.s_lookup_value_valid({firewall_tcpport_table_0lookup_p_0_value_valid}),
	.s_lookup_value_data({firewall_tcpport_table_0lookup_p_0_value_data}),
	.s_lookup_value_ready({firewall_tcpport_table_0lookup_p_0_value_ready}),
	//update port 
	.s_update_req_index({firewall_tcpport_table_0update_p_0_req_index}),
	.s_update_req_index_valid({firewall_tcpport_table_0update_p_0_req_index_valid}),
	.s_update_req_index_ready({firewall_tcpport_table_0update_p_0_req_index_ready}),
	.s_update_req_data({firewall_tcpport_table_0update_p_0_req_data}),
	.s_update_req_data_valid({firewall_tcpport_table_0update_p_0_req_data_valid}),
	.s_update_req_data_ready({firewall_tcpport_table_0update_p_0_req_data_ready})
);

//Table lookup port wire def 
 wire [32-1:0] firewall_tcpport_table_0lookup_p_0_req_index;
 wire  firewall_tcpport_table_0lookup_p_0_req_valid;
 wire  firewall_tcpport_table_0lookup_p_0_req_ready;
 wire  firewall_tcpport_table_0lookup_p_0_value_valid;
 wire  firewall_tcpport_table_0lookup_p_0_value_ready;
 wire [160-1:0] firewall_tcpport_table_0lookup_p_0_value_data;

//Table update port wire def 
 wire [32-1:0] firewall_tcpport_table_0update_p_0_req_index;
 wire  firewall_tcpport_table_0update_p_0_req_index_valid;
 wire  firewall_tcpport_table_0update_p_0_req_index_ready;
 wire [160-1:0] firewall_tcpport_table_0update_p_0_req_data;
 wire  firewall_tcpport_table_0update_p_0_req_data_valid;
 wire  firewall_tcpport_table_0update_p_0_req_data_ready;

atom_CAM#(
)flow_tracker_table_2(
	 .clk(clk), 
	 .rst(rst) ,
	//lookup port 
	.s_lookup_req_index({flow_tracker_table_2lookup_p_0_req_index}),
	.s_lookup_req_valid({flow_tracker_table_2lookup_p_0_req_valid}),
	.s_lookup_req_ready({flow_tracker_table_2lookup_p_0_req_ready}),
	.s_lookup_value_valid({flow_tracker_table_2lookup_p_0_value_valid}),
	.s_lookup_value_data({flow_tracker_table_2lookup_p_0_value_data}),
	.s_lookup_value_ready({flow_tracker_table_2lookup_p_0_value_ready}),
	//update port 
	.s_update_req_index({flow_tracker_table_2update_p_0_req_index}),
	.s_update_req_index_valid({flow_tracker_table_2update_p_0_req_index_valid}),
	.s_update_req_index_ready({flow_tracker_table_2update_p_0_req_index_ready}),
	.s_update_req_data({flow_tracker_table_2update_p_0_req_data}),
	.s_update_req_data_valid({flow_tracker_table_2update_p_0_req_data_valid}),
	.s_update_req_data_ready({flow_tracker_table_2update_p_0_req_data_ready})
);

//Table lookup port wire def 
 wire [32-1:0] flow_tracker_table_2lookup_p_0_req_index;
 wire  flow_tracker_table_2lookup_p_0_req_valid;
 wire  flow_tracker_table_2lookup_p_0_req_ready;
 wire  flow_tracker_table_2lookup_p_0_value_valid;
 wire  flow_tracker_table_2lookup_p_0_value_ready;
 wire [64-1:0] flow_tracker_table_2lookup_p_0_value_data;

//Table update port wire def 
 wire [32-1:0] flow_tracker_table_2update_p_0_req_index;
 wire  flow_tracker_table_2update_p_0_req_index_valid;
 wire  flow_tracker_table_2update_p_0_req_index_ready;
 wire [64-1:0] flow_tracker_table_2update_p_0_req_data;
 wire  flow_tracker_table_2update_p_0_req_data_valid;
 wire  flow_tracker_table_2update_p_0_req_data_ready;

atom_CAM#(
)ip_tracker_table_4(
	 .clk(clk), 
	 .rst(rst) ,
	//lookup port 
	.s_lookup_req_index({ip_tracker_table_4lookup_p_0_req_index}),
	.s_lookup_req_valid({ip_tracker_table_4lookup_p_0_req_valid}),
	.s_lookup_req_ready({ip_tracker_table_4lookup_p_0_req_ready}),
	.s_lookup_value_valid({ip_tracker_table_4lookup_p_0_value_valid}),
	.s_lookup_value_data({ip_tracker_table_4lookup_p_0_value_data}),
	.s_lookup_value_ready({ip_tracker_table_4lookup_p_0_value_ready}),
	//update port 
	.s_update_req_index({ip_tracker_table_4update_p_0_req_index}),
	.s_update_req_index_valid({ip_tracker_table_4update_p_0_req_index_valid}),
	.s_update_req_index_ready({ip_tracker_table_4update_p_0_req_index_ready}),
	.s_update_req_data({ip_tracker_table_4update_p_0_req_data}),
	.s_update_req_data_valid({ip_tracker_table_4update_p_0_req_data_valid}),
	.s_update_req_data_ready({ip_tracker_table_4update_p_0_req_data_ready})
);

//Table lookup port wire def 
 wire [32-1:0] ip_tracker_table_4lookup_p_0_req_index;
 wire  ip_tracker_table_4lookup_p_0_req_valid;
 wire  ip_tracker_table_4lookup_p_0_req_ready;
 wire  ip_tracker_table_4lookup_p_0_value_valid;
 wire  ip_tracker_table_4lookup_p_0_value_ready;
 wire [96-1:0] ip_tracker_table_4lookup_p_0_value_data;

//Table update port wire def 
 wire [32-1:0] ip_tracker_table_4update_p_0_req_index;
 wire  ip_tracker_table_4update_p_0_req_index_valid;
 wire  ip_tracker_table_4update_p_0_req_index_ready;
 wire [96-1:0] ip_tracker_table_4update_p_0_req_data;
 wire  ip_tracker_table_4update_p_0_req_data_valid;
 wire  ip_tracker_table_4update_p_0_req_data_ready;

atom_CAM#(
)lb_fwd_table_7(
	 .clk(clk), 
	 .rst(rst) ,
	//lookup port 
	.s_lookup_req_index({lb_fwd_table_7lookup_p_0_req_index}),
	.s_lookup_req_valid({lb_fwd_table_7lookup_p_0_req_valid}),
	.s_lookup_req_ready({lb_fwd_table_7lookup_p_0_req_ready}),
	.s_lookup_value_valid({lb_fwd_table_7lookup_p_0_value_valid}),
	.s_lookup_value_data({lb_fwd_table_7lookup_p_0_value_data}),
	.s_lookup_value_ready({lb_fwd_table_7lookup_p_0_value_ready}),
	//update port 
	.s_update_req_index({lb_fwd_table_7update_p_0_req_index}),
	.s_update_req_index_valid({lb_fwd_table_7update_p_0_req_index_valid}),
	.s_update_req_index_ready({lb_fwd_table_7update_p_0_req_index_ready}),
	.s_update_req_data({lb_fwd_table_7update_p_0_req_data}),
	.s_update_req_data_valid({lb_fwd_table_7update_p_0_req_data_valid}),
	.s_update_req_data_ready({lb_fwd_table_7update_p_0_req_data_ready})
);

//Table lookup port wire def 
 wire [32-1:0] lb_fwd_table_7lookup_p_0_req_index;
 wire  lb_fwd_table_7lookup_p_0_req_valid;
 wire  lb_fwd_table_7lookup_p_0_req_ready;
 wire  lb_fwd_table_7lookup_p_0_value_valid;
 wire  lb_fwd_table_7lookup_p_0_value_ready;
 wire [160-1:0] lb_fwd_table_7lookup_p_0_value_data;

//Table update port wire def 
 wire [32-1:0] lb_fwd_table_7update_p_0_req_index;
 wire  lb_fwd_table_7update_p_0_req_index_valid;
 wire  lb_fwd_table_7update_p_0_req_index_ready;
 wire [160-1:0] lb_fwd_table_7update_p_0_req_data;
 wire  lb_fwd_table_7update_p_0_req_data_valid;
 wire  lb_fwd_table_7update_p_0_req_data_ready;

atom_CAM#(
)lb_table_6(
	 .clk(clk), 
	 .rst(rst) ,
	//lookup port 
	.s_lookup_req_index({lb_table_6lookup_p_0_req_index}),
	.s_lookup_req_valid({lb_table_6lookup_p_0_req_valid}),
	.s_lookup_req_ready({lb_table_6lookup_p_0_req_ready}),
	.s_lookup_value_valid({lb_table_6lookup_p_0_value_valid}),
	.s_lookup_value_data({lb_table_6lookup_p_0_value_data}),
	.s_lookup_value_ready({lb_table_6lookup_p_0_value_ready}),
	//update port 
	.s_update_req_index({lb_table_6update_p_0_req_index}),
	.s_update_req_index_valid({lb_table_6update_p_0_req_index_valid}),
	.s_update_req_index_ready({lb_table_6update_p_0_req_index_ready}),
	.s_update_req_data({lb_table_6update_p_0_req_data}),
	.s_update_req_data_valid({lb_table_6update_p_0_req_data_valid}),
	.s_update_req_data_ready({lb_table_6update_p_0_req_data_ready})
);

//Table lookup port wire def 
 wire [16-1:0] lb_table_6lookup_p_0_req_index;
 wire  lb_table_6lookup_p_0_req_valid;
 wire  lb_table_6lookup_p_0_req_ready;
 wire  lb_table_6lookup_p_0_value_valid;
 wire  lb_table_6lookup_p_0_value_ready;
 wire [320-1:0] lb_table_6lookup_p_0_value_data;

//Table update port wire def 
 wire [16-1:0] lb_table_6update_p_0_req_index;
 wire  lb_table_6update_p_0_req_index_valid;
 wire  lb_table_6update_p_0_req_index_ready;
 wire [320-1:0] lb_table_6update_p_0_req_data;
 wire  lb_table_6update_p_0_req_data_valid;
 wire  lb_table_6update_p_0_req_data_ready;

atom_CAM#(
)priority_table_1(
	 .clk(clk), 
	 .rst(rst) ,
	//lookup port 
	.s_lookup_req_index({priority_table_1lookup_p_0_req_index}),
	.s_lookup_req_valid({priority_table_1lookup_p_0_req_valid}),
	.s_lookup_req_ready({priority_table_1lookup_p_0_req_ready}),
	.s_lookup_value_valid({priority_table_1lookup_p_0_value_valid}),
	.s_lookup_value_data({priority_table_1lookup_p_0_value_data}),
	.s_lookup_value_ready({priority_table_1lookup_p_0_value_ready}),
	//update port 
	.s_update_req_index({priority_table_1update_p_0_req_index}),
	.s_update_req_index_valid({priority_table_1update_p_0_req_index_valid}),
	.s_update_req_index_ready({priority_table_1update_p_0_req_index_ready}),
	.s_update_req_data({priority_table_1update_p_0_req_data}),
	.s_update_req_data_valid({priority_table_1update_p_0_req_data_valid}),
	.s_update_req_data_ready({priority_table_1update_p_0_req_data_ready})
);

//Table lookup port wire def 
 wire [32-1:0] priority_table_1lookup_p_0_req_index;
 wire  priority_table_1lookup_p_0_req_valid;
 wire  priority_table_1lookup_p_0_req_ready;
 wire  priority_table_1lookup_p_0_value_valid;
 wire  priority_table_1lookup_p_0_value_ready;
 wire [64-1:0] priority_table_1lookup_p_0_value_data;

//Table update port wire def 
 wire [32-1:0] priority_table_1update_p_0_req_index;
 wire  priority_table_1update_p_0_req_index_valid;
 wire  priority_table_1update_p_0_req_index_ready;
 wire [64-1:0] priority_table_1update_p_0_req_data;
 wire  priority_table_1update_p_0_req_data_valid;
 wire  priority_table_1update_p_0_req_data_ready;

atom_CAM#(
)tcp_tracker_table_5(
	 .clk(clk), 
	 .rst(rst) ,
	//lookup port 
	.s_lookup_req_index({tcp_tracker_table_5lookup_p_0_req_index}),
	.s_lookup_req_valid({tcp_tracker_table_5lookup_p_0_req_valid}),
	.s_lookup_req_ready({tcp_tracker_table_5lookup_p_0_req_ready}),
	.s_lookup_value_valid({tcp_tracker_table_5lookup_p_0_value_valid}),
	.s_lookup_value_data({tcp_tracker_table_5lookup_p_0_value_data}),
	.s_lookup_value_ready({tcp_tracker_table_5lookup_p_0_value_ready}),
	//update port 
	.s_update_req_index({tcp_tracker_table_5update_p_0_req_index}),
	.s_update_req_index_valid({tcp_tracker_table_5update_p_0_req_index_valid}),
	.s_update_req_index_ready({tcp_tracker_table_5update_p_0_req_index_ready}),
	.s_update_req_data({tcp_tracker_table_5update_p_0_req_data}),
	.s_update_req_data_valid({tcp_tracker_table_5update_p_0_req_data_valid}),
	.s_update_req_data_ready({tcp_tracker_table_5update_p_0_req_data_ready})
);

//Table lookup port wire def 
 wire [32-1:0] tcp_tracker_table_5lookup_p_0_req_index;
 wire  tcp_tracker_table_5lookup_p_0_req_valid;
 wire  tcp_tracker_table_5lookup_p_0_req_ready;
 wire  tcp_tracker_table_5lookup_p_0_value_valid;
 wire  tcp_tracker_table_5lookup_p_0_value_ready;
 wire [96-1:0] tcp_tracker_table_5lookup_p_0_value_data;

//Table update port wire def 
 wire [32-1:0] tcp_tracker_table_5update_p_0_req_index;
 wire  tcp_tracker_table_5update_p_0_req_index_valid;
 wire  tcp_tracker_table_5update_p_0_req_index_ready;
 wire [96-1:0] tcp_tracker_table_5update_p_0_req_data;
 wire  tcp_tracker_table_5update_p_0_req_data_valid;
 wire  tcp_tracker_table_5update_p_0_req_data_ready;

//
 wire [512-1:0] NET_RECV_0_r0_tdata;
 wire [64-1:0] NET_RECV_0_r0_tkeep;
 wire  NET_RECV_0_r0_tvalid;
 wire  NET_RECV_0_r0_tready;
 wire  NET_RECV_0_r0_tlast;

//
 wire [32-1:0] outport_8_0_r0_tdata;
 wire  outport_8_0_r0_tvalid;
 wire  outport_8_0_r0_tready;

//
 wire [32-1:0] outport_8_1_r0_tdata;
 wire  outport_8_1_r0_tvalid;
 wire  outport_8_1_r0_tready;

//
 wire [32-1:0] outport_8_2_r0_tdata;
 wire  outport_8_2_r0_tvalid;
 wire  outport_8_2_r0_tready;

//
 wire [32-1:0] outport_8_3_r0_tdata;
 wire  outport_8_3_r0_tvalid;
 wire  outport_8_3_r0_tready;

//
 wire [32-1:0] outport_8_4_r0_tdata;
 wire  outport_8_4_r0_tvalid;
 wire  outport_8_4_r0_tready;

//
 wire [32-1:0] outport_8_5_r0_tdata;
 wire  outport_8_5_r0_tvalid;
 wire  outport_8_5_r0_tready;

//
 wire [32-1:0] outport_8_6_r0_tdata;
 wire  outport_8_6_r0_tvalid;
 wire  outport_8_6_r0_tready;

//
 wire [160-1:0] outport_8_7_r0_tdata;
 wire  outport_8_7_r0_tvalid;
 wire  outport_8_7_r0_tready;

//
 wire [512-1:0] outport_8_8_r0_tdata;
 wire [64-1:0] outport_8_8_r0_tkeep;
 wire  outport_8_8_r0_tvalid;
 wire  outport_8_8_r0_tready;
 wire  outport_8_8_r0_tlast;

//
 wire [32-1:0] outport_8_9_r0_tdata;
 wire  outport_8_9_r0_tvalid;
 wire  outport_8_9_r0_tready;

__handler_NET_RECV_process_packet#(
)__handler_NET_RECV_process_packet_351(
	 .clk(clk), 
	 .rst(rst) ,
	//
	.NET_RECV_0_tdata({NET_RECV_0_r0_tdata}),
	.NET_RECV_0_tkeep({NET_RECV_0_r0_tkeep}),
	.NET_RECV_0_tlast({NET_RECV_0_r0_tlast}),
	.NET_RECV_0_tvalid({NET_RECV_0_r0_tvalid}),
	.NET_RECV_0_tready({NET_RECV_0_r0_tready}),
	//
	.outport_8_0_tdata({outport_8_0_r0_tdata}),
	.outport_8_0_tvalid({outport_8_0_r0_tvalid}),
	.outport_8_0_tready({outport_8_0_r0_tready}),
	//
	.outport_8_1_tdata({outport_8_1_r0_tdata}),
	.outport_8_1_tvalid({outport_8_1_r0_tvalid}),
	.outport_8_1_tready({outport_8_1_r0_tready}),
	//
	.outport_8_2_tdata({outport_8_2_r0_tdata}),
	.outport_8_2_tvalid({outport_8_2_r0_tvalid}),
	.outport_8_2_tready({outport_8_2_r0_tready}),
	//
	.outport_8_3_tdata({outport_8_3_r0_tdata}),
	.outport_8_3_tvalid({outport_8_3_r0_tvalid}),
	.outport_8_3_tready({outport_8_3_r0_tready}),
	//
	.outport_8_4_tdata({outport_8_4_r0_tdata}),
	.outport_8_4_tvalid({outport_8_4_r0_tvalid}),
	.outport_8_4_tready({outport_8_4_r0_tready}),
	//
	.outport_8_5_tdata({outport_8_5_r0_tdata}),
	.outport_8_5_tvalid({outport_8_5_r0_tvalid}),
	.outport_8_5_tready({outport_8_5_r0_tready}),
	//
	.outport_8_6_tdata({outport_8_6_r0_tdata}),
	.outport_8_6_tvalid({outport_8_6_r0_tvalid}),
	.outport_8_6_tready({outport_8_6_r0_tready}),
	//
	.outport_8_7_tdata({outport_8_7_r0_tdata}),
	.outport_8_7_tvalid({outport_8_7_r0_tvalid}),
	.outport_8_7_tready({outport_8_7_r0_tready}),
	//
	.outport_8_8_tdata({outport_8_8_r0_tdata}),
	.outport_8_8_tkeep({outport_8_8_r0_tkeep}),
	.outport_8_8_tlast({outport_8_8_r0_tlast}),
	.outport_8_8_tvalid({outport_8_8_r0_tvalid}),
	.outport_8_8_tready({outport_8_8_r0_tready}),
	//
	.outport_8_9_tdata({outport_8_9_r0_tdata}),
	.outport_8_9_tvalid({outport_8_9_r0_tvalid}),
	.outport_8_9_tready({outport_8_9_r0_tready})
);

//
 wire [32-1:0] arg_99_r0_tdata;
 wire  arg_99_r0_tvalid;
 wire  arg_99_r0_tready;

//
 wire [32-1:0] arg_100_r0_tdata;
 wire  arg_100_r0_tvalid;
 wire  arg_100_r0_tready;

//
 wire [32-1:0] arg_101_r0_tdata;
 wire  arg_101_r0_tvalid;
 wire  arg_101_r0_tready;

//
 wire [32-1:0] arg_102_r0_tdata;
 wire  arg_102_r0_tvalid;
 wire  arg_102_r0_tready;

//
 wire [32-1:0] arg_103_r0_tdata;
 wire  arg_103_r0_tvalid;
 wire  arg_103_r0_tready;

//
 wire [32-1:0] arg_104_r0_tdata;
 wire  arg_104_r0_tvalid;
 wire  arg_104_r0_tready;

//
 wire [32-1:0] arg_105_r0_tdata;
 wire  arg_105_r0_tvalid;
 wire  arg_105_r0_tready;

//
 wire [160-1:0] arg_106_r0_tdata;
 wire  arg_106_r0_tvalid;
 wire  arg_106_r0_tready;

//
 wire [512-1:0] arg_107_r0_tdata;
 wire [64-1:0] arg_107_r0_tkeep;
 wire  arg_107_r0_tvalid;
 wire  arg_107_r0_tready;
 wire  arg_107_r0_tlast;

//
 wire [32-1:0] arg_108_r0_tdata;
 wire  arg_108_r0_tvalid;
 wire  arg_108_r0_tready;

//
 wire [32-1:0] outport_109_0_r0_tdata;
 wire  outport_109_0_r0_tvalid;
 wire  outport_109_0_r0_tready;

//
 wire [512-1:0] outport_109_1_r0_tdata;
 wire [64-1:0] outport_109_1_r0_tkeep;
 wire  outport_109_1_r0_tvalid;
 wire  outport_109_1_r0_tready;
 wire  outport_109_1_r0_tlast;

//
 wire [32-1:0] outport_109_2_r0_tdata;
 wire  outport_109_2_r0_tvalid;
 wire  outport_109_2_r0_tready;

//
 wire [32-1:0] outport_109_3_r0_tdata;
 wire  outport_109_3_r0_tvalid;
 wire  outport_109_3_r0_tready;

//
 wire [32-1:0] outport_109_4_r0_tdata;
 wire  outport_109_4_r0_tvalid;
 wire  outport_109_4_r0_tready;

//
 wire [32-1:0] outport_109_5_r0_tdata;
 wire  outport_109_5_r0_tvalid;
 wire  outport_109_5_r0_tready;

//
 wire [32-1:0] outport_109_6_r0_tdata;
 wire  outport_109_6_r0_tvalid;
 wire  outport_109_6_r0_tready;

//
 wire [32-1:0] outport_109_7_r0_tdata;
 wire  outport_109_7_r0_tvalid;
 wire  outport_109_7_r0_tready;

//
 wire [160-1:0] outport_109_8_r0_tdata;
 wire  outport_109_8_r0_tvalid;
 wire  outport_109_8_r0_tready;

__handler_NET_RECV_1_process_packet#(
)__handler_NET_RECV_1_process_packet_352(
	 .clk(clk), 
	 .rst(rst) ,
	//
	.arg_99_tdata({arg_99_r0_tdata}),
	.arg_99_tvalid({arg_99_r0_tvalid}),
	.arg_99_tready({arg_99_r0_tready}),
	//
	.arg_100_tdata({arg_100_r0_tdata}),
	.arg_100_tvalid({arg_100_r0_tvalid}),
	.arg_100_tready({arg_100_r0_tready}),
	//
	.arg_101_tdata({arg_101_r0_tdata}),
	.arg_101_tvalid({arg_101_r0_tvalid}),
	.arg_101_tready({arg_101_r0_tready}),
	//
	.arg_102_tdata({arg_102_r0_tdata}),
	.arg_102_tvalid({arg_102_r0_tvalid}),
	.arg_102_tready({arg_102_r0_tready}),
	//
	.arg_103_tdata({arg_103_r0_tdata}),
	.arg_103_tvalid({arg_103_r0_tvalid}),
	.arg_103_tready({arg_103_r0_tready}),
	//
	.arg_104_tdata({arg_104_r0_tdata}),
	.arg_104_tvalid({arg_104_r0_tvalid}),
	.arg_104_tready({arg_104_r0_tready}),
	//
	.arg_105_tdata({arg_105_r0_tdata}),
	.arg_105_tvalid({arg_105_r0_tvalid}),
	.arg_105_tready({arg_105_r0_tready}),
	//
	.arg_106_tdata({arg_106_r0_tdata}),
	.arg_106_tvalid({arg_106_r0_tvalid}),
	.arg_106_tready({arg_106_r0_tready}),
	//
	.arg_107_tdata({arg_107_r0_tdata}),
	.arg_107_tkeep({arg_107_r0_tkeep}),
	.arg_107_tlast({arg_107_r0_tlast}),
	.arg_107_tvalid({arg_107_r0_tvalid}),
	.arg_107_tready({arg_107_r0_tready}),
	//
	.arg_108_tdata({arg_108_r0_tdata}),
	.arg_108_tvalid({arg_108_r0_tvalid}),
	.arg_108_tready({arg_108_r0_tready}),
	//
	.outport_109_0_tdata({outport_109_0_r0_tdata}),
	.outport_109_0_tvalid({outport_109_0_r0_tvalid}),
	.outport_109_0_tready({outport_109_0_r0_tready}),
	//
	.outport_109_1_tdata({outport_109_1_r0_tdata}),
	.outport_109_1_tkeep({outport_109_1_r0_tkeep}),
	.outport_109_1_tlast({outport_109_1_r0_tlast}),
	.outport_109_1_tvalid({outport_109_1_r0_tvalid}),
	.outport_109_1_tready({outport_109_1_r0_tready}),
	//
	.outport_109_2_tdata({outport_109_2_r0_tdata}),
	.outport_109_2_tvalid({outport_109_2_r0_tvalid}),
	.outport_109_2_tready({outport_109_2_r0_tready}),
	//
	.outport_109_3_tdata({outport_109_3_r0_tdata}),
	.outport_109_3_tvalid({outport_109_3_r0_tvalid}),
	.outport_109_3_tready({outport_109_3_r0_tready}),
	//
	.outport_109_4_tdata({outport_109_4_r0_tdata}),
	.outport_109_4_tvalid({outport_109_4_r0_tvalid}),
	.outport_109_4_tready({outport_109_4_r0_tready}),
	//
	.outport_109_5_tdata({outport_109_5_r0_tdata}),
	.outport_109_5_tvalid({outport_109_5_r0_tvalid}),
	.outport_109_5_tready({outport_109_5_r0_tready}),
	//
	.outport_109_6_tdata({outport_109_6_r0_tdata}),
	.outport_109_6_tvalid({outport_109_6_r0_tvalid}),
	.outport_109_6_tready({outport_109_6_r0_tready}),
	//
	.outport_109_7_tdata({outport_109_7_r0_tdata}),
	.outport_109_7_tvalid({outport_109_7_r0_tvalid}),
	.outport_109_7_tready({outport_109_7_r0_tready}),
	//
	.outport_109_8_tdata({outport_109_8_r0_tdata}),
	.outport_109_8_tvalid({outport_109_8_r0_tvalid}),
	.outport_109_8_tready({outport_109_8_r0_tready})
);

//
 wire [32-1:0] arg_137_r0_tdata;
 wire  arg_137_r0_tvalid;
 wire  arg_137_r0_tready;

//
 wire [512-1:0] arg_138_r0_tdata;
 wire [64-1:0] arg_138_r0_tkeep;
 wire  arg_138_r0_tvalid;
 wire  arg_138_r0_tready;
 wire  arg_138_r0_tlast;

//
 wire [32-1:0] arg_139_r0_tdata;
 wire  arg_139_r0_tvalid;
 wire  arg_139_r0_tready;

//
 wire [32-1:0] arg_140_r0_tdata;
 wire  arg_140_r0_tvalid;
 wire  arg_140_r0_tready;

//
 wire [32-1:0] arg_141_r0_tdata;
 wire  arg_141_r0_tvalid;
 wire  arg_141_r0_tready;

//
 wire [32-1:0] arg_142_r0_tdata;
 wire  arg_142_r0_tvalid;
 wire  arg_142_r0_tready;

//
 wire [32-1:0] arg_143_r0_tdata;
 wire  arg_143_r0_tvalid;
 wire  arg_143_r0_tready;

//
 wire [32-1:0] arg_144_r0_tdata;
 wire  arg_144_r0_tvalid;
 wire  arg_144_r0_tready;

//
 wire [160-1:0] arg_145_r0_tdata;
 wire  arg_145_r0_tvalid;
 wire  arg_145_r0_tready;

//
 wire [32-1:0] outport_146_0_r0_tdata;
 wire  outport_146_0_r0_tvalid;
 wire  outport_146_0_r0_tready;

//
 wire [32-1:0] outport_146_1_r0_tdata;
 wire  outport_146_1_r0_tvalid;
 wire  outport_146_1_r0_tready;

//
 wire [32-1:0] outport_146_2_r0_tdata;
 wire  outport_146_2_r0_tvalid;
 wire  outport_146_2_r0_tready;

//
 wire [32-1:0] outport_146_3_r0_tdata;
 wire  outport_146_3_r0_tvalid;
 wire  outport_146_3_r0_tready;

//
 wire [32-1:0] outport_146_4_r0_tdata;
 wire  outport_146_4_r0_tvalid;
 wire  outport_146_4_r0_tready;

//
 wire [512-1:0] outport_146_5_r0_tdata;
 wire [64-1:0] outport_146_5_r0_tkeep;
 wire  outport_146_5_r0_tvalid;
 wire  outport_146_5_r0_tready;
 wire  outport_146_5_r0_tlast;

//
 wire [160-1:0] outport_146_6_r0_tdata;
 wire  outport_146_6_r0_tvalid;
 wire  outport_146_6_r0_tready;

//
 wire [32-1:0] outport_146_7_r0_tdata;
 wire  outport_146_7_r0_tvalid;
 wire  outport_146_7_r0_tready;

//
 wire [224-1:0] outport_146_8_r0_tdata;
 wire  outport_146_8_r0_tvalid;
 wire  outport_146_8_r0_tready;

__handler_NET_RECV_2_process_packet#(
)__handler_NET_RECV_2_process_packet_353(
	 .clk(clk), 
	 .rst(rst) ,
	//
	.arg_137_tdata({arg_137_r0_tdata}),
	.arg_137_tvalid({arg_137_r0_tvalid}),
	.arg_137_tready({arg_137_r0_tready}),
	//
	.arg_138_tdata({arg_138_r0_tdata}),
	.arg_138_tkeep({arg_138_r0_tkeep}),
	.arg_138_tlast({arg_138_r0_tlast}),
	.arg_138_tvalid({arg_138_r0_tvalid}),
	.arg_138_tready({arg_138_r0_tready}),
	//
	.arg_139_tdata({arg_139_r0_tdata}),
	.arg_139_tvalid({arg_139_r0_tvalid}),
	.arg_139_tready({arg_139_r0_tready}),
	//
	.arg_140_tdata({arg_140_r0_tdata}),
	.arg_140_tvalid({arg_140_r0_tvalid}),
	.arg_140_tready({arg_140_r0_tready}),
	//
	.arg_141_tdata({arg_141_r0_tdata}),
	.arg_141_tvalid({arg_141_r0_tvalid}),
	.arg_141_tready({arg_141_r0_tready}),
	//
	.arg_142_tdata({arg_142_r0_tdata}),
	.arg_142_tvalid({arg_142_r0_tvalid}),
	.arg_142_tready({arg_142_r0_tready}),
	//
	.arg_143_tdata({arg_143_r0_tdata}),
	.arg_143_tvalid({arg_143_r0_tvalid}),
	.arg_143_tready({arg_143_r0_tready}),
	//
	.arg_144_tdata({arg_144_r0_tdata}),
	.arg_144_tvalid({arg_144_r0_tvalid}),
	.arg_144_tready({arg_144_r0_tready}),
	//
	.arg_145_tdata({arg_145_r0_tdata}),
	.arg_145_tvalid({arg_145_r0_tvalid}),
	.arg_145_tready({arg_145_r0_tready}),
	//
	.outport_146_0_tdata({outport_146_0_r0_tdata}),
	.outport_146_0_tvalid({outport_146_0_r0_tvalid}),
	.outport_146_0_tready({outport_146_0_r0_tready}),
	//
	.outport_146_1_tdata({outport_146_1_r0_tdata}),
	.outport_146_1_tvalid({outport_146_1_r0_tvalid}),
	.outport_146_1_tready({outport_146_1_r0_tready}),
	//
	.outport_146_2_tdata({outport_146_2_r0_tdata}),
	.outport_146_2_tvalid({outport_146_2_r0_tvalid}),
	.outport_146_2_tready({outport_146_2_r0_tready}),
	//
	.outport_146_3_tdata({outport_146_3_r0_tdata}),
	.outport_146_3_tvalid({outport_146_3_r0_tvalid}),
	.outport_146_3_tready({outport_146_3_r0_tready}),
	//
	.outport_146_4_tdata({outport_146_4_r0_tdata}),
	.outport_146_4_tvalid({outport_146_4_r0_tvalid}),
	.outport_146_4_tready({outport_146_4_r0_tready}),
	//
	.outport_146_5_tdata({outport_146_5_r0_tdata}),
	.outport_146_5_tkeep({outport_146_5_r0_tkeep}),
	.outport_146_5_tlast({outport_146_5_r0_tlast}),
	.outport_146_5_tvalid({outport_146_5_r0_tvalid}),
	.outport_146_5_tready({outport_146_5_r0_tready}),
	//
	.outport_146_6_tdata({outport_146_6_r0_tdata}),
	.outport_146_6_tvalid({outport_146_6_r0_tvalid}),
	.outport_146_6_tready({outport_146_6_r0_tready}),
	//
	.outport_146_7_tdata({outport_146_7_r0_tdata}),
	.outport_146_7_tvalid({outport_146_7_r0_tvalid}),
	.outport_146_7_tready({outport_146_7_r0_tready}),
	//
	.outport_146_8_tdata({outport_146_8_r0_tdata}),
	.outport_146_8_tvalid({outport_146_8_r0_tvalid}),
	.outport_146_8_tready({outport_146_8_r0_tready})
);

//
 wire [32-1:0] arg_162_r0_tdata;
 wire  arg_162_r0_tvalid;
 wire  arg_162_r0_tready;

//
 wire [32-1:0] arg_163_r0_tdata;
 wire  arg_163_r0_tvalid;
 wire  arg_163_r0_tready;

//
 wire [32-1:0] arg_164_r0_tdata;
 wire  arg_164_r0_tvalid;
 wire  arg_164_r0_tready;

//
 wire [32-1:0] arg_165_r0_tdata;
 wire  arg_165_r0_tvalid;
 wire  arg_165_r0_tready;

//
 wire [32-1:0] arg_166_r0_tdata;
 wire  arg_166_r0_tvalid;
 wire  arg_166_r0_tready;

//
 wire [512-1:0] arg_167_r0_tdata;
 wire [64-1:0] arg_167_r0_tkeep;
 wire  arg_167_r0_tvalid;
 wire  arg_167_r0_tready;
 wire  arg_167_r0_tlast;

//
 wire [160-1:0] arg_168_r0_tdata;
 wire  arg_168_r0_tvalid;
 wire  arg_168_r0_tready;

//
 wire [32-1:0] arg_169_r0_tdata;
 wire  arg_169_r0_tvalid;
 wire  arg_169_r0_tready;

//
 wire [224-1:0] arg_170_r0_tdata;
 wire  arg_170_r0_tvalid;
 wire  arg_170_r0_tready;

//
 wire [512-1:0] NET_SEND_0_r0_tdata;
 wire [64-1:0] NET_SEND_0_r0_tkeep;
 wire  NET_SEND_0_r0_tvalid;
 wire  NET_SEND_0_r0_tready;
 wire  NET_SEND_0_r0_tlast;

__handler_NET_RECV_3_process_packet#(
)__handler_NET_RECV_3_process_packet_354(
	 .clk(clk), 
	 .rst(rst) ,
	//
	.arg_162_tdata({arg_162_r0_tdata}),
	.arg_162_tvalid({arg_162_r0_tvalid}),
	.arg_162_tready({arg_162_r0_tready}),
	//
	.arg_163_tdata({arg_163_r0_tdata}),
	.arg_163_tvalid({arg_163_r0_tvalid}),
	.arg_163_tready({arg_163_r0_tready}),
	//
	.arg_164_tdata({arg_164_r0_tdata}),
	.arg_164_tvalid({arg_164_r0_tvalid}),
	.arg_164_tready({arg_164_r0_tready}),
	//
	.arg_165_tdata({arg_165_r0_tdata}),
	.arg_165_tvalid({arg_165_r0_tvalid}),
	.arg_165_tready({arg_165_r0_tready}),
	//
	.arg_166_tdata({arg_166_r0_tdata}),
	.arg_166_tvalid({arg_166_r0_tvalid}),
	.arg_166_tready({arg_166_r0_tready}),
	//
	.arg_167_tdata({arg_167_r0_tdata}),
	.arg_167_tkeep({arg_167_r0_tkeep}),
	.arg_167_tlast({arg_167_r0_tlast}),
	.arg_167_tvalid({arg_167_r0_tvalid}),
	.arg_167_tready({arg_167_r0_tready}),
	//
	.arg_168_tdata({arg_168_r0_tdata}),
	.arg_168_tvalid({arg_168_r0_tvalid}),
	.arg_168_tready({arg_168_r0_tready}),
	//
	.arg_169_tdata({arg_169_r0_tdata}),
	.arg_169_tvalid({arg_169_r0_tvalid}),
	.arg_169_tready({arg_169_r0_tready}),
	//
	.arg_170_tdata({arg_170_r0_tdata}),
	.arg_170_tvalid({arg_170_r0_tvalid}),
	.arg_170_tready({arg_170_r0_tready}),
	//
	.NET_SEND_0_tdata({NET_SEND_0_r0_tdata}),
	.NET_SEND_0_tkeep({NET_SEND_0_r0_tkeep}),
	.NET_SEND_0_tlast({NET_SEND_0_r0_tlast}),
	.NET_SEND_0_tvalid({NET_SEND_0_r0_tvalid}),
	.NET_SEND_0_tready({NET_SEND_0_r0_tready})
);

//
 wire [32-1:0] in_0_arg_99_tdata;
 wire  in_0_arg_99_tvalid;
 wire  in_0_arg_99_tready;

//
 wire [32-1:0] in_0_arg_100_tdata;
 wire  in_0_arg_100_tvalid;
 wire  in_0_arg_100_tready;

//
 wire [32-1:0] in_0_arg_101_tdata;
 wire  in_0_arg_101_tvalid;
 wire  in_0_arg_101_tready;

//
 wire [32-1:0] in_0_arg_102_tdata;
 wire  in_0_arg_102_tvalid;
 wire  in_0_arg_102_tready;

//
 wire [32-1:0] in_0_arg_103_tdata;
 wire  in_0_arg_103_tvalid;
 wire  in_0_arg_103_tready;

//
 wire [32-1:0] in_0_arg_104_tdata;
 wire  in_0_arg_104_tvalid;
 wire  in_0_arg_104_tready;

//
 wire [32-1:0] in_0_arg_105_tdata;
 wire  in_0_arg_105_tvalid;
 wire  in_0_arg_105_tready;

//
 wire [160-1:0] in_0_arg_106_tdata;
 wire  in_0_arg_106_tvalid;
 wire  in_0_arg_106_tready;

//
 wire [512-1:0] in_0_arg_107_tdata;
 wire [64-1:0] in_0_arg_107_tkeep;
 wire  in_0_arg_107_tvalid;
 wire  in_0_arg_107_tready;
 wire  in_0_arg_107_tlast;

//
 wire [32-1:0] in_0_arg_108_tdata;
 wire  in_0_arg_108_tvalid;
 wire  in_0_arg_108_tready;

//
 wire [32-1:0] out_0_arg_99_tdata;
 wire  out_0_arg_99_tvalid;
 wire  out_0_arg_99_tready;

//
 wire [32-1:0] out_0_arg_100_tdata;
 wire  out_0_arg_100_tvalid;
 wire  out_0_arg_100_tready;

//
 wire [32-1:0] out_0_arg_101_tdata;
 wire  out_0_arg_101_tvalid;
 wire  out_0_arg_101_tready;

//
 wire [32-1:0] out_0_arg_102_tdata;
 wire  out_0_arg_102_tvalid;
 wire  out_0_arg_102_tready;

//
 wire [32-1:0] out_0_arg_103_tdata;
 wire  out_0_arg_103_tvalid;
 wire  out_0_arg_103_tready;

//
 wire [32-1:0] out_0_arg_104_tdata;
 wire  out_0_arg_104_tvalid;
 wire  out_0_arg_104_tready;

//
 wire [32-1:0] out_0_arg_105_tdata;
 wire  out_0_arg_105_tvalid;
 wire  out_0_arg_105_tready;

//
 wire [160-1:0] out_0_arg_106_tdata;
 wire  out_0_arg_106_tvalid;
 wire  out_0_arg_106_tready;

//
 wire [512-1:0] out_0_arg_107_tdata;
 wire [64-1:0] out_0_arg_107_tkeep;
 wire  out_0_arg_107_tvalid;
 wire  out_0_arg_107_tready;
 wire  out_0_arg_107_tlast;

//
 wire [32-1:0] out_0_arg_108_tdata;
 wire  out_0_arg_108_tvalid;
 wire  out_0_arg_108_tready;

__controller_NET_RECV_1#(
)__controller_NET_RECV_1_355(
	 .clk(clk), 
	 .rst(rst) ,
	//
	.in_0_arg_99_tdata({in_0_arg_99_tdata}),
	.in_0_arg_99_tvalid({in_0_arg_99_tvalid}),
	.in_0_arg_99_tready({in_0_arg_99_tready}),
	//
	.in_0_arg_100_tdata({in_0_arg_100_tdata}),
	.in_0_arg_100_tvalid({in_0_arg_100_tvalid}),
	.in_0_arg_100_tready({in_0_arg_100_tready}),
	//
	.in_0_arg_101_tdata({in_0_arg_101_tdata}),
	.in_0_arg_101_tvalid({in_0_arg_101_tvalid}),
	.in_0_arg_101_tready({in_0_arg_101_tready}),
	//
	.in_0_arg_102_tdata({in_0_arg_102_tdata}),
	.in_0_arg_102_tvalid({in_0_arg_102_tvalid}),
	.in_0_arg_102_tready({in_0_arg_102_tready}),
	//
	.in_0_arg_103_tdata({in_0_arg_103_tdata}),
	.in_0_arg_103_tvalid({in_0_arg_103_tvalid}),
	.in_0_arg_103_tready({in_0_arg_103_tready}),
	//
	.in_0_arg_104_tdata({in_0_arg_104_tdata}),
	.in_0_arg_104_tvalid({in_0_arg_104_tvalid}),
	.in_0_arg_104_tready({in_0_arg_104_tready}),
	//
	.in_0_arg_105_tdata({in_0_arg_105_tdata}),
	.in_0_arg_105_tvalid({in_0_arg_105_tvalid}),
	.in_0_arg_105_tready({in_0_arg_105_tready}),
	//
	.in_0_arg_106_tdata({in_0_arg_106_tdata}),
	.in_0_arg_106_tvalid({in_0_arg_106_tvalid}),
	.in_0_arg_106_tready({in_0_arg_106_tready}),
	//
	.in_0_arg_107_tdata({in_0_arg_107_tdata}),
	.in_0_arg_107_tkeep({in_0_arg_107_tkeep}),
	.in_0_arg_107_tlast({in_0_arg_107_tlast}),
	.in_0_arg_107_tvalid({in_0_arg_107_tvalid}),
	.in_0_arg_107_tready({in_0_arg_107_tready}),
	//
	.in_0_arg_108_tdata({in_0_arg_108_tdata}),
	.in_0_arg_108_tvalid({in_0_arg_108_tvalid}),
	.in_0_arg_108_tready({in_0_arg_108_tready}),
	//
	.out_0_arg_99_tdata({out_0_arg_99_tdata}),
	.out_0_arg_99_tvalid({out_0_arg_99_tvalid}),
	.out_0_arg_99_tready({out_0_arg_99_tready}),
	//
	.out_0_arg_100_tdata({out_0_arg_100_tdata}),
	.out_0_arg_100_tvalid({out_0_arg_100_tvalid}),
	.out_0_arg_100_tready({out_0_arg_100_tready}),
	//
	.out_0_arg_101_tdata({out_0_arg_101_tdata}),
	.out_0_arg_101_tvalid({out_0_arg_101_tvalid}),
	.out_0_arg_101_tready({out_0_arg_101_tready}),
	//
	.out_0_arg_102_tdata({out_0_arg_102_tdata}),
	.out_0_arg_102_tvalid({out_0_arg_102_tvalid}),
	.out_0_arg_102_tready({out_0_arg_102_tready}),
	//
	.out_0_arg_103_tdata({out_0_arg_103_tdata}),
	.out_0_arg_103_tvalid({out_0_arg_103_tvalid}),
	.out_0_arg_103_tready({out_0_arg_103_tready}),
	//
	.out_0_arg_104_tdata({out_0_arg_104_tdata}),
	.out_0_arg_104_tvalid({out_0_arg_104_tvalid}),
	.out_0_arg_104_tready({out_0_arg_104_tready}),
	//
	.out_0_arg_105_tdata({out_0_arg_105_tdata}),
	.out_0_arg_105_tvalid({out_0_arg_105_tvalid}),
	.out_0_arg_105_tready({out_0_arg_105_tready}),
	//
	.out_0_arg_106_tdata({out_0_arg_106_tdata}),
	.out_0_arg_106_tvalid({out_0_arg_106_tvalid}),
	.out_0_arg_106_tready({out_0_arg_106_tready}),
	//
	.out_0_arg_107_tdata({out_0_arg_107_tdata}),
	.out_0_arg_107_tkeep({out_0_arg_107_tkeep}),
	.out_0_arg_107_tlast({out_0_arg_107_tlast}),
	.out_0_arg_107_tvalid({out_0_arg_107_tvalid}),
	.out_0_arg_107_tready({out_0_arg_107_tready}),
	//
	.out_0_arg_108_tdata({out_0_arg_108_tdata}),
	.out_0_arg_108_tvalid({out_0_arg_108_tvalid}),
	.out_0_arg_108_tready({out_0_arg_108_tready})
);

//
 wire [32-1:0] in_0_arg_137_tdata;
 wire  in_0_arg_137_tvalid;
 wire  in_0_arg_137_tready;

//
 wire [512-1:0] in_0_arg_138_tdata;
 wire [64-1:0] in_0_arg_138_tkeep;
 wire  in_0_arg_138_tvalid;
 wire  in_0_arg_138_tready;
 wire  in_0_arg_138_tlast;

//
 wire [32-1:0] in_0_arg_139_tdata;
 wire  in_0_arg_139_tvalid;
 wire  in_0_arg_139_tready;

//
 wire [32-1:0] in_0_arg_140_tdata;
 wire  in_0_arg_140_tvalid;
 wire  in_0_arg_140_tready;

//
 wire [32-1:0] in_0_arg_141_tdata;
 wire  in_0_arg_141_tvalid;
 wire  in_0_arg_141_tready;

//
 wire [32-1:0] in_0_arg_142_tdata;
 wire  in_0_arg_142_tvalid;
 wire  in_0_arg_142_tready;

//
 wire [32-1:0] in_0_arg_143_tdata;
 wire  in_0_arg_143_tvalid;
 wire  in_0_arg_143_tready;

//
 wire [32-1:0] in_0_arg_144_tdata;
 wire  in_0_arg_144_tvalid;
 wire  in_0_arg_144_tready;

//
 wire [160-1:0] in_0_arg_145_tdata;
 wire  in_0_arg_145_tvalid;
 wire  in_0_arg_145_tready;

//
 wire [32-1:0] out_0_arg_137_tdata;
 wire  out_0_arg_137_tvalid;
 wire  out_0_arg_137_tready;

//
 wire [512-1:0] out_0_arg_138_tdata;
 wire [64-1:0] out_0_arg_138_tkeep;
 wire  out_0_arg_138_tvalid;
 wire  out_0_arg_138_tready;
 wire  out_0_arg_138_tlast;

//
 wire [32-1:0] out_0_arg_139_tdata;
 wire  out_0_arg_139_tvalid;
 wire  out_0_arg_139_tready;

//
 wire [32-1:0] out_0_arg_140_tdata;
 wire  out_0_arg_140_tvalid;
 wire  out_0_arg_140_tready;

//
 wire [32-1:0] out_0_arg_141_tdata;
 wire  out_0_arg_141_tvalid;
 wire  out_0_arg_141_tready;

//
 wire [32-1:0] out_0_arg_142_tdata;
 wire  out_0_arg_142_tvalid;
 wire  out_0_arg_142_tready;

//
 wire [32-1:0] out_0_arg_143_tdata;
 wire  out_0_arg_143_tvalid;
 wire  out_0_arg_143_tready;

//
 wire [32-1:0] out_0_arg_144_tdata;
 wire  out_0_arg_144_tvalid;
 wire  out_0_arg_144_tready;

//
 wire [160-1:0] out_0_arg_145_tdata;
 wire  out_0_arg_145_tvalid;
 wire  out_0_arg_145_tready;

__controller_NET_RECV_2#(
)__controller_NET_RECV_2_356(
	 .clk(clk), 
	 .rst(rst) ,
	//
	.in_0_arg_137_tdata({in_0_arg_137_tdata}),
	.in_0_arg_137_tvalid({in_0_arg_137_tvalid}),
	.in_0_arg_137_tready({in_0_arg_137_tready}),
	//
	.in_0_arg_138_tdata({in_0_arg_138_tdata}),
	.in_0_arg_138_tkeep({in_0_arg_138_tkeep}),
	.in_0_arg_138_tlast({in_0_arg_138_tlast}),
	.in_0_arg_138_tvalid({in_0_arg_138_tvalid}),
	.in_0_arg_138_tready({in_0_arg_138_tready}),
	//
	.in_0_arg_139_tdata({in_0_arg_139_tdata}),
	.in_0_arg_139_tvalid({in_0_arg_139_tvalid}),
	.in_0_arg_139_tready({in_0_arg_139_tready}),
	//
	.in_0_arg_140_tdata({in_0_arg_140_tdata}),
	.in_0_arg_140_tvalid({in_0_arg_140_tvalid}),
	.in_0_arg_140_tready({in_0_arg_140_tready}),
	//
	.in_0_arg_141_tdata({in_0_arg_141_tdata}),
	.in_0_arg_141_tvalid({in_0_arg_141_tvalid}),
	.in_0_arg_141_tready({in_0_arg_141_tready}),
	//
	.in_0_arg_142_tdata({in_0_arg_142_tdata}),
	.in_0_arg_142_tvalid({in_0_arg_142_tvalid}),
	.in_0_arg_142_tready({in_0_arg_142_tready}),
	//
	.in_0_arg_143_tdata({in_0_arg_143_tdata}),
	.in_0_arg_143_tvalid({in_0_arg_143_tvalid}),
	.in_0_arg_143_tready({in_0_arg_143_tready}),
	//
	.in_0_arg_144_tdata({in_0_arg_144_tdata}),
	.in_0_arg_144_tvalid({in_0_arg_144_tvalid}),
	.in_0_arg_144_tready({in_0_arg_144_tready}),
	//
	.in_0_arg_145_tdata({in_0_arg_145_tdata}),
	.in_0_arg_145_tvalid({in_0_arg_145_tvalid}),
	.in_0_arg_145_tready({in_0_arg_145_tready}),
	//
	.out_0_arg_137_tdata({out_0_arg_137_tdata}),
	.out_0_arg_137_tvalid({out_0_arg_137_tvalid}),
	.out_0_arg_137_tready({out_0_arg_137_tready}),
	//
	.out_0_arg_138_tdata({out_0_arg_138_tdata}),
	.out_0_arg_138_tkeep({out_0_arg_138_tkeep}),
	.out_0_arg_138_tlast({out_0_arg_138_tlast}),
	.out_0_arg_138_tvalid({out_0_arg_138_tvalid}),
	.out_0_arg_138_tready({out_0_arg_138_tready}),
	//
	.out_0_arg_139_tdata({out_0_arg_139_tdata}),
	.out_0_arg_139_tvalid({out_0_arg_139_tvalid}),
	.out_0_arg_139_tready({out_0_arg_139_tready}),
	//
	.out_0_arg_140_tdata({out_0_arg_140_tdata}),
	.out_0_arg_140_tvalid({out_0_arg_140_tvalid}),
	.out_0_arg_140_tready({out_0_arg_140_tready}),
	//
	.out_0_arg_141_tdata({out_0_arg_141_tdata}),
	.out_0_arg_141_tvalid({out_0_arg_141_tvalid}),
	.out_0_arg_141_tready({out_0_arg_141_tready}),
	//
	.out_0_arg_142_tdata({out_0_arg_142_tdata}),
	.out_0_arg_142_tvalid({out_0_arg_142_tvalid}),
	.out_0_arg_142_tready({out_0_arg_142_tready}),
	//
	.out_0_arg_143_tdata({out_0_arg_143_tdata}),
	.out_0_arg_143_tvalid({out_0_arg_143_tvalid}),
	.out_0_arg_143_tready({out_0_arg_143_tready}),
	//
	.out_0_arg_144_tdata({out_0_arg_144_tdata}),
	.out_0_arg_144_tvalid({out_0_arg_144_tvalid}),
	.out_0_arg_144_tready({out_0_arg_144_tready}),
	//
	.out_0_arg_145_tdata({out_0_arg_145_tdata}),
	.out_0_arg_145_tvalid({out_0_arg_145_tvalid}),
	.out_0_arg_145_tready({out_0_arg_145_tready})
);

//
 wire [32-1:0] in_0_arg_162_tdata;
 wire  in_0_arg_162_tvalid;
 wire  in_0_arg_162_tready;

//
 wire [32-1:0] in_0_arg_163_tdata;
 wire  in_0_arg_163_tvalid;
 wire  in_0_arg_163_tready;

//
 wire [32-1:0] in_0_arg_164_tdata;
 wire  in_0_arg_164_tvalid;
 wire  in_0_arg_164_tready;

//
 wire [32-1:0] in_0_arg_165_tdata;
 wire  in_0_arg_165_tvalid;
 wire  in_0_arg_165_tready;

//
 wire [32-1:0] in_0_arg_166_tdata;
 wire  in_0_arg_166_tvalid;
 wire  in_0_arg_166_tready;

//
 wire [512-1:0] in_0_arg_167_tdata;
 wire [64-1:0] in_0_arg_167_tkeep;
 wire  in_0_arg_167_tvalid;
 wire  in_0_arg_167_tready;
 wire  in_0_arg_167_tlast;

//
 wire [160-1:0] in_0_arg_168_tdata;
 wire  in_0_arg_168_tvalid;
 wire  in_0_arg_168_tready;

//
 wire [32-1:0] in_0_arg_169_tdata;
 wire  in_0_arg_169_tvalid;
 wire  in_0_arg_169_tready;

//
 wire [224-1:0] in_0_arg_170_tdata;
 wire  in_0_arg_170_tvalid;
 wire  in_0_arg_170_tready;

//
 wire [32-1:0] out_0_arg_162_tdata;
 wire  out_0_arg_162_tvalid;
 wire  out_0_arg_162_tready;

//
 wire [32-1:0] out_0_arg_163_tdata;
 wire  out_0_arg_163_tvalid;
 wire  out_0_arg_163_tready;

//
 wire [32-1:0] out_0_arg_164_tdata;
 wire  out_0_arg_164_tvalid;
 wire  out_0_arg_164_tready;

//
 wire [32-1:0] out_0_arg_165_tdata;
 wire  out_0_arg_165_tvalid;
 wire  out_0_arg_165_tready;

//
 wire [32-1:0] out_0_arg_166_tdata;
 wire  out_0_arg_166_tvalid;
 wire  out_0_arg_166_tready;

//
 wire [512-1:0] out_0_arg_167_tdata;
 wire [64-1:0] out_0_arg_167_tkeep;
 wire  out_0_arg_167_tvalid;
 wire  out_0_arg_167_tready;
 wire  out_0_arg_167_tlast;

//
 wire [160-1:0] out_0_arg_168_tdata;
 wire  out_0_arg_168_tvalid;
 wire  out_0_arg_168_tready;

//
 wire [32-1:0] out_0_arg_169_tdata;
 wire  out_0_arg_169_tvalid;
 wire  out_0_arg_169_tready;

//
 wire [224-1:0] out_0_arg_170_tdata;
 wire  out_0_arg_170_tvalid;
 wire  out_0_arg_170_tready;

__controller_NET_RECV_3#(
)__controller_NET_RECV_3_357(
	 .clk(clk), 
	 .rst(rst) ,
	//
	.in_0_arg_162_tdata({in_0_arg_162_tdata}),
	.in_0_arg_162_tvalid({in_0_arg_162_tvalid}),
	.in_0_arg_162_tready({in_0_arg_162_tready}),
	//
	.in_0_arg_163_tdata({in_0_arg_163_tdata}),
	.in_0_arg_163_tvalid({in_0_arg_163_tvalid}),
	.in_0_arg_163_tready({in_0_arg_163_tready}),
	//
	.in_0_arg_164_tdata({in_0_arg_164_tdata}),
	.in_0_arg_164_tvalid({in_0_arg_164_tvalid}),
	.in_0_arg_164_tready({in_0_arg_164_tready}),
	//
	.in_0_arg_165_tdata({in_0_arg_165_tdata}),
	.in_0_arg_165_tvalid({in_0_arg_165_tvalid}),
	.in_0_arg_165_tready({in_0_arg_165_tready}),
	//
	.in_0_arg_166_tdata({in_0_arg_166_tdata}),
	.in_0_arg_166_tvalid({in_0_arg_166_tvalid}),
	.in_0_arg_166_tready({in_0_arg_166_tready}),
	//
	.in_0_arg_167_tdata({in_0_arg_167_tdata}),
	.in_0_arg_167_tkeep({in_0_arg_167_tkeep}),
	.in_0_arg_167_tlast({in_0_arg_167_tlast}),
	.in_0_arg_167_tvalid({in_0_arg_167_tvalid}),
	.in_0_arg_167_tready({in_0_arg_167_tready}),
	//
	.in_0_arg_168_tdata({in_0_arg_168_tdata}),
	.in_0_arg_168_tvalid({in_0_arg_168_tvalid}),
	.in_0_arg_168_tready({in_0_arg_168_tready}),
	//
	.in_0_arg_169_tdata({in_0_arg_169_tdata}),
	.in_0_arg_169_tvalid({in_0_arg_169_tvalid}),
	.in_0_arg_169_tready({in_0_arg_169_tready}),
	//
	.in_0_arg_170_tdata({in_0_arg_170_tdata}),
	.in_0_arg_170_tvalid({in_0_arg_170_tvalid}),
	.in_0_arg_170_tready({in_0_arg_170_tready}),
	//
	.out_0_arg_162_tdata({out_0_arg_162_tdata}),
	.out_0_arg_162_tvalid({out_0_arg_162_tvalid}),
	.out_0_arg_162_tready({out_0_arg_162_tready}),
	//
	.out_0_arg_163_tdata({out_0_arg_163_tdata}),
	.out_0_arg_163_tvalid({out_0_arg_163_tvalid}),
	.out_0_arg_163_tready({out_0_arg_163_tready}),
	//
	.out_0_arg_164_tdata({out_0_arg_164_tdata}),
	.out_0_arg_164_tvalid({out_0_arg_164_tvalid}),
	.out_0_arg_164_tready({out_0_arg_164_tready}),
	//
	.out_0_arg_165_tdata({out_0_arg_165_tdata}),
	.out_0_arg_165_tvalid({out_0_arg_165_tvalid}),
	.out_0_arg_165_tready({out_0_arg_165_tready}),
	//
	.out_0_arg_166_tdata({out_0_arg_166_tdata}),
	.out_0_arg_166_tvalid({out_0_arg_166_tvalid}),
	.out_0_arg_166_tready({out_0_arg_166_tready}),
	//
	.out_0_arg_167_tdata({out_0_arg_167_tdata}),
	.out_0_arg_167_tkeep({out_0_arg_167_tkeep}),
	.out_0_arg_167_tlast({out_0_arg_167_tlast}),
	.out_0_arg_167_tvalid({out_0_arg_167_tvalid}),
	.out_0_arg_167_tready({out_0_arg_167_tready}),
	//
	.out_0_arg_168_tdata({out_0_arg_168_tdata}),
	.out_0_arg_168_tvalid({out_0_arg_168_tvalid}),
	.out_0_arg_168_tready({out_0_arg_168_tready}),
	//
	.out_0_arg_169_tdata({out_0_arg_169_tdata}),
	.out_0_arg_169_tvalid({out_0_arg_169_tvalid}),
	.out_0_arg_169_tready({out_0_arg_169_tready}),
	//
	.out_0_arg_170_tdata({out_0_arg_170_tdata}),
	.out_0_arg_170_tvalid({out_0_arg_170_tvalid}),
	.out_0_arg_170_tready({out_0_arg_170_tready})
);

 assign in_0_arg_99_tdata = outport_8_0_r0_tdata;
 assign in_0_arg_99_tvalid = outport_8_0_r0_tvalid;
 assign outport_8_0_r0_tready = in_0_arg_99_tready;

 assign in_0_arg_100_tdata = outport_8_1_r0_tdata;
 assign in_0_arg_100_tvalid = outport_8_1_r0_tvalid;
 assign outport_8_1_r0_tready = in_0_arg_100_tready;

 assign in_0_arg_101_tdata = outport_8_2_r0_tdata;
 assign in_0_arg_101_tvalid = outport_8_2_r0_tvalid;
 assign outport_8_2_r0_tready = in_0_arg_101_tready;

 assign in_0_arg_102_tdata = outport_8_3_r0_tdata;
 assign in_0_arg_102_tvalid = outport_8_3_r0_tvalid;
 assign outport_8_3_r0_tready = in_0_arg_102_tready;

 assign in_0_arg_103_tdata = outport_8_4_r0_tdata;
 assign in_0_arg_103_tvalid = outport_8_4_r0_tvalid;
 assign outport_8_4_r0_tready = in_0_arg_103_tready;

 assign in_0_arg_104_tdata = outport_8_5_r0_tdata;
 assign in_0_arg_104_tvalid = outport_8_5_r0_tvalid;
 assign outport_8_5_r0_tready = in_0_arg_104_tready;

 assign in_0_arg_105_tdata = outport_8_6_r0_tdata;
 assign in_0_arg_105_tvalid = outport_8_6_r0_tvalid;
 assign outport_8_6_r0_tready = in_0_arg_105_tready;

 assign in_0_arg_106_tdata = outport_8_7_r0_tdata;
 assign in_0_arg_106_tvalid = outport_8_7_r0_tvalid;
 assign outport_8_7_r0_tready = in_0_arg_106_tready;

 assign in_0_arg_107_tdata = outport_8_8_r0_tdata;
 assign in_0_arg_107_tvalid = outport_8_8_r0_tvalid;
 assign outport_8_8_r0_tready = in_0_arg_107_tready;
 assign in_0_arg_107_tkeep = outport_8_8_r0_tkeep;
 assign in_0_arg_107_tlast = outport_8_8_r0_tlast;

 assign in_0_arg_108_tdata = outport_8_9_r0_tdata;
 assign in_0_arg_108_tvalid = outport_8_9_r0_tvalid;
 assign outport_8_9_r0_tready = in_0_arg_108_tready;

 assign arg_99_r0_tdata = out_0_arg_99_tdata;
 assign arg_99_r0_tvalid = out_0_arg_99_tvalid;
 assign out_0_arg_99_tready = arg_99_r0_tready;

 assign arg_100_r0_tdata = out_0_arg_100_tdata;
 assign arg_100_r0_tvalid = out_0_arg_100_tvalid;
 assign out_0_arg_100_tready = arg_100_r0_tready;

 assign arg_101_r0_tdata = out_0_arg_101_tdata;
 assign arg_101_r0_tvalid = out_0_arg_101_tvalid;
 assign out_0_arg_101_tready = arg_101_r0_tready;

 assign arg_102_r0_tdata = out_0_arg_102_tdata;
 assign arg_102_r0_tvalid = out_0_arg_102_tvalid;
 assign out_0_arg_102_tready = arg_102_r0_tready;

 assign arg_103_r0_tdata = out_0_arg_103_tdata;
 assign arg_103_r0_tvalid = out_0_arg_103_tvalid;
 assign out_0_arg_103_tready = arg_103_r0_tready;

 assign arg_104_r0_tdata = out_0_arg_104_tdata;
 assign arg_104_r0_tvalid = out_0_arg_104_tvalid;
 assign out_0_arg_104_tready = arg_104_r0_tready;

 assign arg_105_r0_tdata = out_0_arg_105_tdata;
 assign arg_105_r0_tvalid = out_0_arg_105_tvalid;
 assign out_0_arg_105_tready = arg_105_r0_tready;

 assign arg_106_r0_tdata = out_0_arg_106_tdata;
 assign arg_106_r0_tvalid = out_0_arg_106_tvalid;
 assign out_0_arg_106_tready = arg_106_r0_tready;

 assign arg_107_r0_tdata = out_0_arg_107_tdata;
 assign arg_107_r0_tvalid = out_0_arg_107_tvalid;
 assign out_0_arg_107_tready = arg_107_r0_tready;
 assign arg_107_r0_tkeep = out_0_arg_107_tkeep;
 assign arg_107_r0_tlast = out_0_arg_107_tlast;

 assign arg_108_r0_tdata = out_0_arg_108_tdata;
 assign arg_108_r0_tvalid = out_0_arg_108_tvalid;
 assign out_0_arg_108_tready = arg_108_r0_tready;

 assign in_0_arg_137_tdata = outport_109_0_r0_tdata;
 assign in_0_arg_137_tvalid = outport_109_0_r0_tvalid;
 assign outport_109_0_r0_tready = in_0_arg_137_tready;

 assign in_0_arg_138_tdata = outport_109_1_r0_tdata;
 assign in_0_arg_138_tvalid = outport_109_1_r0_tvalid;
 assign outport_109_1_r0_tready = in_0_arg_138_tready;
 assign in_0_arg_138_tkeep = outport_109_1_r0_tkeep;
 assign in_0_arg_138_tlast = outport_109_1_r0_tlast;

 assign in_0_arg_139_tdata = outport_109_2_r0_tdata;
 assign in_0_arg_139_tvalid = outport_109_2_r0_tvalid;
 assign outport_109_2_r0_tready = in_0_arg_139_tready;

 assign in_0_arg_140_tdata = outport_109_3_r0_tdata;
 assign in_0_arg_140_tvalid = outport_109_3_r0_tvalid;
 assign outport_109_3_r0_tready = in_0_arg_140_tready;

 assign in_0_arg_141_tdata = outport_109_4_r0_tdata;
 assign in_0_arg_141_tvalid = outport_109_4_r0_tvalid;
 assign outport_109_4_r0_tready = in_0_arg_141_tready;

 assign in_0_arg_142_tdata = outport_109_5_r0_tdata;
 assign in_0_arg_142_tvalid = outport_109_5_r0_tvalid;
 assign outport_109_5_r0_tready = in_0_arg_142_tready;

 assign in_0_arg_143_tdata = outport_109_6_r0_tdata;
 assign in_0_arg_143_tvalid = outport_109_6_r0_tvalid;
 assign outport_109_6_r0_tready = in_0_arg_143_tready;

 assign in_0_arg_144_tdata = outport_109_7_r0_tdata;
 assign in_0_arg_144_tvalid = outport_109_7_r0_tvalid;
 assign outport_109_7_r0_tready = in_0_arg_144_tready;

 assign in_0_arg_145_tdata = outport_109_8_r0_tdata;
 assign in_0_arg_145_tvalid = outport_109_8_r0_tvalid;
 assign outport_109_8_r0_tready = in_0_arg_145_tready;

 assign arg_137_r0_tdata = out_0_arg_137_tdata;
 assign arg_137_r0_tvalid = out_0_arg_137_tvalid;
 assign out_0_arg_137_tready = arg_137_r0_tready;

 assign arg_138_r0_tdata = out_0_arg_138_tdata;
 assign arg_138_r0_tvalid = out_0_arg_138_tvalid;
 assign out_0_arg_138_tready = arg_138_r0_tready;
 assign arg_138_r0_tkeep = out_0_arg_138_tkeep;
 assign arg_138_r0_tlast = out_0_arg_138_tlast;

 assign arg_139_r0_tdata = out_0_arg_139_tdata;
 assign arg_139_r0_tvalid = out_0_arg_139_tvalid;
 assign out_0_arg_139_tready = arg_139_r0_tready;

 assign arg_140_r0_tdata = out_0_arg_140_tdata;
 assign arg_140_r0_tvalid = out_0_arg_140_tvalid;
 assign out_0_arg_140_tready = arg_140_r0_tready;

 assign arg_141_r0_tdata = out_0_arg_141_tdata;
 assign arg_141_r0_tvalid = out_0_arg_141_tvalid;
 assign out_0_arg_141_tready = arg_141_r0_tready;

 assign arg_142_r0_tdata = out_0_arg_142_tdata;
 assign arg_142_r0_tvalid = out_0_arg_142_tvalid;
 assign out_0_arg_142_tready = arg_142_r0_tready;

 assign arg_143_r0_tdata = out_0_arg_143_tdata;
 assign arg_143_r0_tvalid = out_0_arg_143_tvalid;
 assign out_0_arg_143_tready = arg_143_r0_tready;

 assign arg_144_r0_tdata = out_0_arg_144_tdata;
 assign arg_144_r0_tvalid = out_0_arg_144_tvalid;
 assign out_0_arg_144_tready = arg_144_r0_tready;

 assign arg_145_r0_tdata = out_0_arg_145_tdata;
 assign arg_145_r0_tvalid = out_0_arg_145_tvalid;
 assign out_0_arg_145_tready = arg_145_r0_tready;

 assign in_0_arg_162_tdata = outport_146_0_r0_tdata;
 assign in_0_arg_162_tvalid = outport_146_0_r0_tvalid;
 assign outport_146_0_r0_tready = in_0_arg_162_tready;

 assign in_0_arg_163_tdata = outport_146_1_r0_tdata;
 assign in_0_arg_163_tvalid = outport_146_1_r0_tvalid;
 assign outport_146_1_r0_tready = in_0_arg_163_tready;

 assign in_0_arg_164_tdata = outport_146_2_r0_tdata;
 assign in_0_arg_164_tvalid = outport_146_2_r0_tvalid;
 assign outport_146_2_r0_tready = in_0_arg_164_tready;

 assign in_0_arg_165_tdata = outport_146_3_r0_tdata;
 assign in_0_arg_165_tvalid = outport_146_3_r0_tvalid;
 assign outport_146_3_r0_tready = in_0_arg_165_tready;

 assign in_0_arg_166_tdata = outport_146_4_r0_tdata;
 assign in_0_arg_166_tvalid = outport_146_4_r0_tvalid;
 assign outport_146_4_r0_tready = in_0_arg_166_tready;

 assign in_0_arg_167_tdata = outport_146_5_r0_tdata;
 assign in_0_arg_167_tvalid = outport_146_5_r0_tvalid;
 assign outport_146_5_r0_tready = in_0_arg_167_tready;
 assign in_0_arg_167_tkeep = outport_146_5_r0_tkeep;
 assign in_0_arg_167_tlast = outport_146_5_r0_tlast;

 assign in_0_arg_168_tdata = outport_146_6_r0_tdata;
 assign in_0_arg_168_tvalid = outport_146_6_r0_tvalid;
 assign outport_146_6_r0_tready = in_0_arg_168_tready;

 assign in_0_arg_169_tdata = outport_146_7_r0_tdata;
 assign in_0_arg_169_tvalid = outport_146_7_r0_tvalid;
 assign outport_146_7_r0_tready = in_0_arg_169_tready;

 assign in_0_arg_170_tdata = outport_146_8_r0_tdata;
 assign in_0_arg_170_tvalid = outport_146_8_r0_tvalid;
 assign outport_146_8_r0_tready = in_0_arg_170_tready;

 assign arg_162_r0_tdata = out_0_arg_162_tdata;
 assign arg_162_r0_tvalid = out_0_arg_162_tvalid;
 assign out_0_arg_162_tready = arg_162_r0_tready;

 assign arg_163_r0_tdata = out_0_arg_163_tdata;
 assign arg_163_r0_tvalid = out_0_arg_163_tvalid;
 assign out_0_arg_163_tready = arg_163_r0_tready;

 assign arg_164_r0_tdata = out_0_arg_164_tdata;
 assign arg_164_r0_tvalid = out_0_arg_164_tvalid;
 assign out_0_arg_164_tready = arg_164_r0_tready;

 assign arg_165_r0_tdata = out_0_arg_165_tdata;
 assign arg_165_r0_tvalid = out_0_arg_165_tvalid;
 assign out_0_arg_165_tready = arg_165_r0_tready;

 assign arg_166_r0_tdata = out_0_arg_166_tdata;
 assign arg_166_r0_tvalid = out_0_arg_166_tvalid;
 assign out_0_arg_166_tready = arg_166_r0_tready;

 assign arg_167_r0_tdata = out_0_arg_167_tdata;
 assign arg_167_r0_tvalid = out_0_arg_167_tvalid;
 assign out_0_arg_167_tready = arg_167_r0_tready;
 assign arg_167_r0_tkeep = out_0_arg_167_tkeep;
 assign arg_167_r0_tlast = out_0_arg_167_tlast;

 assign arg_168_r0_tdata = out_0_arg_168_tdata;
 assign arg_168_r0_tvalid = out_0_arg_168_tvalid;
 assign out_0_arg_168_tready = arg_168_r0_tready;

 assign arg_169_r0_tdata = out_0_arg_169_tdata;
 assign arg_169_r0_tvalid = out_0_arg_169_tvalid;
 assign out_0_arg_169_tready = arg_169_r0_tready;

 assign arg_170_r0_tdata = out_0_arg_170_tdata;
 assign arg_170_r0_tvalid = out_0_arg_170_tvalid;
 assign out_0_arg_170_tready = arg_170_r0_tready;

 assign NET_RECV_0_r0_tdata = NET_RECV_0_tdata;
 assign NET_RECV_0_r0_tvalid = NET_RECV_0_tvalid;
 assign NET_RECV_0_tready = NET_RECV_0_r0_tready;
 assign NET_RECV_0_r0_tkeep = NET_RECV_0_tkeep;
 assign NET_RECV_0_r0_tlast = NET_RECV_0_tlast;

 assign NET_SEND_0_tdata = NET_SEND_0_r0_tdata;
 assign NET_SEND_0_tvalid = NET_SEND_0_r0_tvalid;
 assign NET_SEND_0_r0_tready = NET_SEND_0_tready;
 assign NET_SEND_0_tkeep = NET_SEND_0_r0_tkeep;
 assign NET_SEND_0_tlast = NET_SEND_0_r0_tlast;


endmodule
